//Testbench Recorrido Izquierda a Derecha

`timescale 1 ns / 1 ps

module izq_der_tb;

reg [2:0] a, b;
wire w, z;